`timescale 1ns / 1ns 

module tb;

parameter N = 8;

reg [N-1:0] A1, B1;
wire [N-1:0] sum1;

reg [N-1:0] A2, B2;
wire [N-1:0] sum2;

reg [N-1:0] A3, B3;
wire [N-1:0] sum3;

wire [N-1:0] sumActual;
assign sumActual = A1 + B1;

nBitRcpa1 #(.N(N)) nBitRcpa1Inst(
    .A(A1),
    .B(B1),
    .sum(sum1)
);

nBitRcpa2 #(.N(N)) nBitRcpa2Inst(
    .A(A2),
    .B(B2),
    .sum(sum2)
);

nBitRcpa3 #(.N(N)) nBitRcpa3Inst(
    .A(A3),
    .B(B3),
    .sum(sum3)
);


initial begin
    $dumpfile("output.vcd");
    $dumpvars(0, tb);

    // A = 4'b0011; B = 4'b0110; #10;
    // A = 8'b01011110; B = 8'b00110010; #10;
    // A = 1'b1; B = 1'b1; #10; 

	A1 = 8'b00110000; B1 = 8'b00000101; 
	A2 = 8'b00110000; B2 = 8'b00000101;
	A3 = 8'b00110000; B3 = 8'b00000101; #10;
	A1 = 8'b01000111; B1 = 8'b01110000; 
	A2 = 8'b01000111; B2 = 8'b01110000;
	A3 = 8'b01000111; B3 = 8'b01110000; #10;
	A1 = 8'b01000000; B1 = 8'b01110111; 
	A2 = 8'b01000000; B2 = 8'b01110111;
	A3 = 8'b01000000; B3 = 8'b01110111; #10;
	A1 = 8'b00010100; B1 = 8'b01000010; 
	A2 = 8'b00010100; B2 = 8'b01000010;
	A3 = 8'b00010100; B3 = 8'b01000010; #10;
	A1 = 8'b01011001; B1 = 8'b00010111; 
	A2 = 8'b01011001; B2 = 8'b00010111;
	A3 = 8'b01011001; B3 = 8'b00010111; #10;
	A1 = 8'b01001101; B1 = 8'b01100010; 
	A2 = 8'b01001101; B2 = 8'b01100010;
	A3 = 8'b01001101; B3 = 8'b01100010; #10;
	A1 = 8'b01000101; B1 = 8'b00011111; 
	A2 = 8'b01000101; B2 = 8'b00011111;
	A3 = 8'b01000101; B3 = 8'b00011111; #10;
	A1 = 8'b01111000; B1 = 8'b00111000; 
	A2 = 8'b01111000; B2 = 8'b00111000;
	A3 = 8'b01111000; B3 = 8'b00111000; #10;
	A1 = 8'b00001001; B1 = 8'b01110011; 
	A2 = 8'b00001001; B2 = 8'b01110011;
	A3 = 8'b00001001; B3 = 8'b01110011; #10;
	A1 = 8'b00110101; B1 = 8'b01111000; 
	A2 = 8'b00110101; B2 = 8'b01111000;
	A3 = 8'b00110101; B3 = 8'b01111000; #10;


    $finish;
end

endmodule
