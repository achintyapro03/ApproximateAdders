`timescale 1ns / 1ns 

module testbenchhybridfa;

parameter N1= 16,N2=16,addOrSub=0;

reg [N1+N2-1:0] A1, B1;
wire [N1+N2-1:0] sum1;
wire cout1;

reg [N1+N2-1:0] A2, B2;
wire [N1+N2:0] sum2;

assign sum2 = A2 + B2;


HybridAdder #(.N1(N1), .N2(N2), .addOrSub(addOrSub)) HybridAdderInst1(
    .A(A1),
    .B(B1),
    .sum(sum1),
    .cout(cout1)
);


initial begin
    $dumpfile("exe/output_hybrid.vcd");
    $dumpvars(0, testbenchhybridfa);
    // Test vectors with delays
    A1 = 32'b 1010111000110010001000011000001; B1 = 32'b 1110001101111101100000001011101; 
	A2 = 32'b 1010111000110010001000011000001; B2 = 32'b 1110001101111101100000001011101; #10;
	A1 = 32'b 1110100111101111111000000101101; B1 = 32'b 1011000000101000101000000000010; 
	A2 = 32'b 1110100111101111111000000101101; B2 = 32'b 1011000000101000101000000000010; #10;
	A1 = 32'b  101000111010000001010011010110; B1 = 32'b  111001100111100111111101111000; 
	A2 = 32'b  101000111010000001010011010110; B2 = 32'b  111001100111100111111101111000; #10;
	A1 = 32'b   10111001000010000000001010000; B1 = 32'b  100111010101101001111101010111; 
	A2 = 32'b   10111001000010000000001010000; B2 = 32'b  100111010101101001111101010111; #10;
	A1 = 32'b 1101001111100000010000000110010; B1 = 32'b      10011001100101010111110010; 
	A2 = 32'b 1101001111100000010000000110010; B2 = 32'b      10011001100101010111110010; #10;
	A1 = 32'b   11011111000111001011011011100; B1 = 32'b   11000000111111010111101101001; 
	A2 = 32'b   11011111000111001011011011100; B2 = 32'b   11000000111111010111101101001; #10;
	A1 = 32'b 1000101011011010011111100001110; B1 = 32'b  111001101111111111011111000000; 
	A2 = 32'b 1000101011011010011111100001110; B2 = 32'b  111001101111111111011111000000; #10;
	A1 = 32'b 1101101011110110000001111001100; B1 = 32'b 1010001010001000011100111110000; 
	A2 = 32'b 1101101011110110000001111001100; B2 = 32'b 1010001010001000011100111110000; #10;
	A1 = 32'b   10110011010101000010111110001; B1 = 32'b 1100110110010100011111111100010; 
	A2 = 32'b   10110011010101000010111110001; B2 = 32'b 1100110110010100011111111100010; #10;
	A1 = 32'b 1100001000111001011100110011001; B1 = 32'b    1101100100101110011100110011; 
	A2 = 32'b 1100001000111001011100110011001; B2 = 32'b    1101100100101110011100110011; #10;
	A1 = 32'b    1100110010010100000110000011; B1 = 32'b 1001110001111111011010111100100; 
	A2 = 32'b    1100110010010100000110000011; B2 = 32'b 1001110001111111011010111100100; #10;
	A1 = 32'b 1011000110010111101011100010101; B1 = 32'b  100011110010110000011000111000; 
	A2 = 32'b 1011000110010111101011100010101; B2 = 32'b  100011110010110000011000111000; #10;
	A1 = 32'b  111110100101001100100010000101; B1 = 32'b 1100001010101001001001000101011; 
	A2 = 32'b  111110100101001100100010000101; B2 = 32'b 1100001010101001001001000101011; #10;
	A1 = 32'b 1010001100010110001110111100111; B1 = 32'b 1100000011110100011001101001100; 
	A2 = 32'b 1010001100010110001110111100111; B2 = 32'b 1100000011110100011001101001100; #10;
	A1 = 32'b  111101001111110101110100100101; B1 = 32'b       1101011000000000010000011; 
	A2 = 32'b  111101001111110101110100100101; B2 = 32'b       1101011000000000010000011; #10;
	A1 = 32'b 1101110001011111010101110010101; B1 = 32'b 1011011000010110111110101100101; 
	A2 = 32'b 1101110001011111010101110010101; B2 = 32'b 1011011000010110111110101100101; #10;
	A1 = 32'b  111110010001001011101111000111; B1 = 32'b 1100110101111001011111011111010; 
	A2 = 32'b  111110010001001011101111000111; B2 = 32'b 1100110101111001011111011111010; #10;
	A1 = 32'b 1101101000101000011110011111001; B1 = 32'b       1011111101010001011011100; 
	A2 = 32'b 1101101000101000011110011111001; B2 = 32'b       1011111101010001011011100; #10;
	A1 = 32'b   10111101111110101111100101110; B1 = 32'b  101110000100001011111011110111; 
	A2 = 32'b   10111101111110101111100101110; B2 = 32'b  101110000100001011111011110111; #10;
	A1 = 32'b  110101101100011100111001011000; B1 = 32'b 1000101001101011111101011000001; 
	A2 = 32'b  110101101100011100111001011000; B2 = 32'b 1000101001101011111101011000001; #10;



    // Finish simulation
    $finish;
end

endmodule
